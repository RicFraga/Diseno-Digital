LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DECO IS
PORT (
	d, clk: IN STD_LOGIC;
	q: OUT STD_LOGIC
);	
END DECO;

ARCHITECTURE ADECO OF DECO IS
BEGIN	
	PROCESS(clk,d)
		BEGIN IF(clk'event and clk = '1')
			THEN
				q <= d;
		END IF;
	END PROCESS;
END ADECO;