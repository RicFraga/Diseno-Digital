module ru ( 
	d0,
	d1,
	d2,
	d3,
	es,
	oper0,
	oper1,
	clk,
	clr,
	q0,
	q1,
	q2,
	q3
	) ;

input  d0;
input  d1;
input  d2;
input  d3;
input  es;
input  oper0;
input  oper1;
input  clk;
input  clr;
inout  q0;
inout  q1;
inout  q2;
inout  q3;
